module timer (
	input clock_25mhz,   // system clock
	input rest_sync,     // system reset
	input [3:0] value,   // initial value
	input start_timer,   // asserted high to start the timer
	output expired       // asserted high when timer ends
	);

	

endmodule

